

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


package wm_package is

constant Data_Width: integer:=32;
    constant shift_param:integer:=16;
  constant  NN_size:integer:=100;
 constant   connection_size:integer:=20;
 constant astro_size:integer:=9;

  type index_array is array (0 to NN_size*connection_size-1) of integer range 0 to 100;------------------ array for saving neuron outputs
 
--constant pre_indx: index_array:=(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,4,4,4,4,4,4,4,4,4,4,4,4,4,4,4,5,5,5,5,5,5,5,5,5,5,5,5,5,5,5,6,6,6,6,6,6,6,6,6,6,6,6,6,6,6,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,8,8,8,8,8,8,8,8,8,8,8,8,8,8,8,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,10,10,10,10,10,10,10,10,10,10,10,10,10,10,10,11,11,11,11,11,11,11,11,11,11,11,11,11,11,11,12,12,12,12,12,12,12,12,12,12,12,12,12,12,12,13,13,13,13,13,13,13,13,13,13,13,13,13,13,13,14,14,14,14,14,14,14,14,14,14,14,14,14,14,14,15,15,15,15,15,15,15,15,15,15,15,15,15,15,15,16,16,16,16,16,16,16,16,16,16,16,16,16,16,16,17,17,17,17,17,17,17,17,17,17,17,17,17,17,17,18,18,18,18,18,18,18,18,18,18,18,18,18,18,18,19,19,19,19,19,19,19,19,19,19,19,19,19,19,19,20,20,20,20,20,20,20,20,20,20,20,20,20,20,20,21,21,21,21,21,21,21,21,21,21,21,21,21,21,21,22,22,22,22,22,22,22,22,22,22,22,22,22,22,22,23,23,23,23,23,23,23,23,23,23,23,23,23,23,23,24,24,24,24,24,24,24,24,24,24,24,24,24,24,24,25,25,25,25,25,25,25,25,25,25,25,25,25,25,25,26,26,26,26,26,26,26,26,26,26,26,26,26,26,26,27,27,27,27,27,27,27,27,27,27,27,27,27,27,27,28,28,28,28,28,28,28,28,28,28,28,28,28,28,28,29,29,29,29,29,29,29,29,29,29,29,29,29,29,29,30,30,30,30,30,30,30,30,30,30,30,30,30,30,30,31,31,31,31,31,31,31,31,31,31,31,31,31,31,31,32,32,32,32,32,32,32,32,32,32,32,32,32,32,32,33,33,33,33,33,33,33,33,33,33,33,33,33,33,33,34,34,34,34,34,34,34,34,34,34,34,34,34,34,34,35,35,35,35,35,35,35,35,35,35,35,35,35,35,35,36,36,36,36,36,36,36,36,36,36,36,36,36,36,36,37,37,37,37,37,37,37,37,37,37,37,37,37,37,37,38,38,38,38,38,38,38,38,38,38,38,38,38,38,38,39,39,39,39,39,39,39,39,39,39,39,39,39,39,39,40,40,40,40,40,40,40,40,40,40,40,40,40,40,40,41,41,41,41,41,41,41,41,41,41,41,41,41,41,41,42,42,42,42,42,42,42,42,42,42,42,42,42,42,42,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43,44,44,44,44,44,44,44,44,44,44,44,44,44,44,44,45,45,45,45,45,45,45,45,45,45,45,45,45,45,45,46,46,46,46,46,46,46,46,46,46,46,46,46,46,46,47,47,47,47,47,47,47,47,47,47,47,47,47,47,47,48,48,48,48,48,48,48,48,48,48,48,48,48,48,48,49,49,49,49,49,49,49,49,49,49,49,49,49,49,49,50,50,50,50,50,50,50,50,50,50,50,50,50,50,50,51,51,51,51,51,51,51,51,51,51,51,51,51,51,51,52,52,52,52,52,52,52,52,52,52,52,52,52,52,52,53,53,53,53,53,53,53,53,53,53,53,53,53,53,53,54,54,54,54,54,54,54,54,54,54,54,54,54,54,54,55,55,55,55,55,55,55,55,55,55,55,55,55,55,55,56,56,56,56,56,56,56,56,56,56,56,56,56,56,56,57,57,57,57,57,57,57,57,57,57,57,57,57,57,57,58,58,58,58,58,58,58,58,58,58,58,58,58,58,58,59,59,59,59,59,59,59,59,59,59,59,59,59,59,59,60,60,60,60,60,60,60,60,60,60,60,60,60,60,60,61,61,61,61,61,61,61,61,61,61,61,61,61,61,61,62,62,62,62,62,62,62,62,62,62,62,62,62,62,62,63,63,63,63,63,63,63,63,63,63,63,63,63,63,63,64,64,64,64,64,64,64,64,64,64,64,64,64,64,64,65,65,65,65,65,65,65,65,65,65,65,65,65,65,65,66,66,66,66,66,66,66,66,66,66,66,66,66,66,66,67,67,67,67,67,67,67,67,67,67,67,67,67,67,67,68,68,68,68,68,68,68,68,68,68,68,68,68,68,68,69,69,69,69,69,69,69,69,69,69,69,69,69,69,69,70,70,70,70,70,70,70,70,70,70,70,70,70,70,70,71,71,71,71,71,71,71,71,71,71,71,71,71,71,71,72,72,72,72,72,72,72,72,72,72,72,72,72,72,72,73,73,73,73,73,73,73,73,73,73,73,73,73,73,73,74,74,74,74,74,74,74,74,74,74,74,74,74,74,74,75,75,75,75,75,75,75,75,75,75,75,75,75,75,75,76,76,76,76,76,76,76,76,76,76,76,76,76,76,76,77,77,77,77,77,77,77,77,77,77,77,77,77,77,77,78,78,78,78,78,78,78,78,78,78,78,78,78,78,78,79,79,79,79,79,79,79,79,79,79,79,79,79,79,79,80,80,80,80,80,80,80,80,80,80,80,80,80,80,80,81,81,81,81,81,81,81,81,81,81,81,81,81,81,81,82,82,82,82,82,82,82,82,82,82,82,82,82,82,82,83,83,83,83,83,83,83,83,83,83,83,83,83,83,83,84,84,84,84,84,84,84,84,84,84,84,84,84,84,84,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,86,86,86,86,86,86,86,86,86,86,86,86,86,86,86,87,87,87,87,87,87,87,87,87,87,87,87,87,87,87,88,88,88,88,88,88,88,88,88,88,88,88,88,88,88,89,89,89,89,89,89,89,89,89,89,89,89,89,89,89,90,90,90,90,90,90,90,90,90,90,90,90,90,90,90,91,91,91,91,91,91,91,91,91,91,91,91,91,91,91,92,92,92,92,92,92,92,92,92,92,92,92,92,92,92,93,93,93,93,93,93,93,93,93,93,93,93,93,93,93,94,94,94,94,94,94,94,94,94,94,94,94,94,94,94,95,95,95,95,95,95,95,95,95,95,95,95,95,95,95,96,96,96,96,96,96,96,96,96,96,96,96,96,96,96,97,97,97,97,97,97,97,97,97,97,97,97,97,97,97,98,98,98,98,98,98,98,98,98,98,98,98,98,98,98,99,99,99,99,99,99,99,99,99,99,99,99,99,99,99,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100);
------------------- post indexes from matlabb
--constant post_indx: index_array:=(11,17,35,2,21,25,3,38,24,12,4,22,31,6,61,41,7,33,13,45,78,62,42,23,80,40,68,5,76,10,42,26,54,1,51,73,3,11,4,22,31,37,35,52,23,93,84,14,43,12,34,45,21,44,6,32,71,56,91,15,4,13,10,26,5,9,11,2,33,21,45,1,24,61,71,34,25,23,8,30,14,27,31,64,60,40,22,58,16,90,8,73,14,82,21,69,5,34,6,3,33,10,2,15,63,11,18,23,54,98,1,62,68,36,45,61,75,48,99,100,66,35,6,23,86,13,14,8,9,38,28,15,84,93,25,87,24,4,16,55,2,7,94,26,19,63,33,39,3,56,15,18,26,9,46,7,39,3,5,27,4,45,1,36,20,96,60,16,84,2,24,25,44,38,14,41,8,11,10,76,37,19,62,47,17,14,18,8,22,48,51,6,70,46,34,4,57,5,9,15,83,27,26,72,49,10,16,3,20,24,9,42,53,48,7,14,57,28,6,18,4,38,62,29,58,3,17,49,34,100,27,43,10,33,37,25,85,19,2,1,44,8,30,7,29,2,57,40,59,10,50,69,19,15,27,58,18,46,24,88,6,63,11,49,4,39,5,37,21,20,4,7,9,50,8,3,29,20,31,19,18,37,30,89,78,46,40,17,5,44,38,74,69,66,27,88,52,36,1,71,25,51,37,41,21,23,1,43,13,14,28,62,53,94,35,32,15,12,65,7,4,2,31,33,52,6,71,24,74,75,11,7,69,23,43,32,22,16,55,24,35,39,1,6,42,45,87,52,2,17,14,33,15,34,82,73,13,61,21,5,95,3,17,25,15,32,35,22,5,21,12,38,14,62,33,49,23,43,2,47,8,96,81,11,52,27,44,72,78,26,75,15,25,36,3,11,44,23,24,37,13,35,10,28,29,7,73,16,4,66,2,17,9,6,53,85,54,26,92,34,16,23,12,27,25,14,90,19,5,97,75,17,31,67,4,32,21,57,6,7,26,38,55,56,35,28,18,58,13,22,5,52,17,29,18,6,8,69,38,15,26,45,2,37,50,30,48,46,14,7,25,59,32,36,19,4,22,49,10,24,39,38,30,28,16,15,63,7,26,6,25,23,4,46,54,67,27,3,8,45,35,57,29,5,50,24,47,94,19,51,17,13,15,5,28,56,88,20,49,58,8,9,12,98,30,35,7,33,68,32,3,29,89,19,87,24,10,93,16,78,20,36,17,27,89,28,29,46,30,50,39,9,14,18,91,12,80,8,98,70,5,52,6,34,69,4,37,26,25,74,10,94,38,19,22,36,30,86,5,89,99,77,55,29,17,9,93,75,23,47,60,26,8,16,69,87,27,40,2,6,51,12,35,23,4,27,43,65,15,52,34,62,2,84,18,11,41,83,22,54,25,44,31,53,97,74,49,32,1,33,31,23,32,21,57,12,51,42,13,43,37,11,7,24,44,72,15,3,5,25,14,92,1,56,33,16,41,52,82,47,31,24,33,43,27,59,77,29,41,7,72,26,13,12,15,3,11,22,21,37,42,88,5,96,32,81,14,25,36,2,44,64,77,14,82,26,45,55,42,32,25,53,35,34,13,19,27,74,22,21,28,43,6,16,41,75,2,4,33,65,33,45,42,75,26,58,35,43,50,40,27,73,98,29,46,23,4,15,10,53,55,59,85,34,87,84,5,61,56,65,49,56,27,21,19,25,4,35,33,17,15,36,6,77,84,28,24,74,79,82,20,66,99,7,16,37,39,94,5,72,26,17,29,59,7,11,18,58,30,28,22,36,78,45,40,37,6,25,24,48,35,68,38,19,67,47,20,74,75,49,95,38,59,9,66,58,41,77,27,24,30,36,13,3,34,5,50,47,17,18,45,2,39,16,52,25,19,15,8,48,56,58,18,39,88,14,19,17,33,30,59,46,28,36,2,38,7,25,40,43,49,5,69,57,27,26,48,79,60,95,51,39,42,82,38,40,60,8,23,29,7,18,26,49,28,31,47,58,80,24,65,10,20,50,67,84,33,9,44,85,33,41,32,1,42,52,58,21,25,15,35,28,66,44,22,34,63,11,71,55,83,62,92,2,36,98,61,49,46,14,14,26,31,42,11,5,12,34,33,24,85,22,51,52,23,81,55,8,29,35,36,41,47,2,79,27,92,9,15,43,23,4,41,30,52,31,37,71,54,44,35,53,32,36,5,72,42,3,25,12,81,49,38,90,26,22,77,16,8,34,24,35,53,94,15,25,42,13,97,62,16,45,36,44,32,43,55,12,57,64,96,37,4,59,54,92,58,26,28,9,64,33,13,69,54,29,47,44,52,25,1,42,79,37,10,51,55,34,94,19,36,39,56,38,45,5,46,67,21,53,25,45,18,33,34,11,80,35,63,30,76,42,98,74,3,4,69,46,38,68,37,53,17,20,24,26,49,65,86,44,35,59,85,47,36,79,98,40,24,16,30,65,7,27,56,8,6,57,38,77,100,46,9,67,26,22,21,39,58,49,48,18,27,56,31,58,40,50,37,46,84,70,49,32,20,28,55,39,59,88,52,69,47,94,30,64,8,10,17,34,49,86,29,59,37,89,98,35,17,40,48,27,38,68,8,15,58,57,30,91,26,100,24,88,34,6,79,70,54,50,50,87,39,6,46,70,38,47,30,60,68,26,17,48,8,79,20,25,43,9,19,100,15,33,49,29,14,66,55,67,52,21,31,64,51,15,34,42,81,45,83,43,11,13,1,48,71,23,44,22,35,61,54,3,33,26,10,12,46,53,8,49,61,22,12,62,32,43,21,53,47,1,2,37,71,82,38,41,80,44,72,56,34,46,35,73,33,25,54,45,44,3,23,55,70,33,17,62,54,94,37,42,27,92,57,14,11,83,77,41,12,2,13,65,35,31,82,46,66,45,34,54,37,43,78,84,45,42,33,47,58,31,4,14,46,28,9,32,74,71,60,24,77,81,64,66,41,59,48,75,77,76,35,55,44,46,38,71,66,93,36,26,51,31,54,33,34,72,56,16,43,42,58,24,20,79,65,53,52,15,75,21,77,45,40,74,78,56,47,13,16,54,70,95,87,28,60,67,100,35,72,53,32,36,27,15,58,43,64,57,50,40,48,27,44,53,58,75,77,49,79,57,94,41,24,45,9,46,37,82,56,80,14,59,36,85,67,13,100,21,58,46,47,65,10,28,82,38,49,26,75,76,68,59,70,64,66,78,41,45,43,40,8,29,74,67,18,57,55,39,48,9,80,47,57,77,29,36,20,79,32,50,46,40,60,38,19,30,59,52,69,27,39,13,58,93,45,55,6,34,46,59,60,70,20,39,40,47,30,49,100,57,10,73,69,15,80,56,48,75,38,37,90,42,87,45,36,41,35,65,31,71,83,63,41,11,33,44,1,61,35,76,32,21,52,78,22,64,37,13,55,65,81,92,16,96,34,62,53,19,93,34,42,59,22,53,62,31,58,55,51,72,18,54,94,56,61,71,63,82,65,24,32,47,8,3,43,75,25,66,56,34,33,43,79,44,52,51,54,6,63,68,98,92,45,13,81,72,31,82,14,5,41,24,55,94,23,87,58,35,74,34,56,42,18,64,47,44,41,62,95,22,14,36,33,88,16,53,59,57,75,52,24,60,91,27,98,87,86,30,28,65,35,25,43,54,66,45,57,44,99,1,63,46,68,47,59,56,37,76,83,75,51,85,93,52,39,64,53,29,66,38,76,46,82,15,55,86,53,94,67,57,26,88,85,18,73,62,47,58,42,50,16,36,48,59,71,68,35,25,50,37,24,75,87,80,67,56,59,90,36,58,46,55,48,42,60,76,38,91,7,30,94,86,53,43,66,65,70,45,37,98,48,60,68,52,51,55,89,67,88,45,50,57,26,49,69,43,28,35,53,39,23,94,36,9,14,84,66,47,48,46,68,58,19,60,49,89,57,99,10,69,13,7,16,47,39,70,9,25,98,67,38,40,79,29,66,88,96,77,57,83,70,93,75,48,68,47,84,28,59,89,40,30,90,58,50,49,65,35,29,52,19,88,78,38,18,51,15,79,5,74,71,51,57,81,90,62,33,77,44,52,1,94,64,48,75,82,36,41,42,84,49,55,24,21,72,78,63,4,63,72,53,73,65,91,41,61,24,20,92,4,33,23,64,43,25,55,32,69,96,42,51,94,79,76,12,58,81,67,74,62,81,64,23,34,94,83,73,82,85,52,33,66,58,45,43,21,56,12,54,78,11,42,48,4,72,68,96,92,66,63,86,67,11,74,54,62,42,65,47,59,24,91,75,34,46,61,84,53,31,73,4,79,50,45,56,10,16,87,54,56,36,85,76,82,66,95,67,39,55,75,61,57,62,77,37,41,2,94,25,53,70,64,97,48,50,91,35,44,70,76,89,86,87,36,97,62,56,48,40,49,18,22,67,65,74,19,46,37,47,24,75,43,69,64,57,55,68,77,83,78,50,68,55,69,77,76,37,43,87,49,19,60,58,39,27,63,98,71,97,6,66,57,75,82,44,45,94,56,99,58,67,54,69,48,88,26,78,11,12,70,79,76,86,63,96,66,38,36,57,30,24,9,75,55,82,50,89,4,59,96,79,21,68,40,58,84,70,66,49,38,88,89,48,6,80,37,67,65,18,77,78,87,30,53,76,29,17,34,60,28,65,59,87,94,69,68,80,34,67,27,100,6,64,4,62,90,98,99,84,29,50,10,79,85,97,30,9,2,62,41,80,91,61,21,82,81,13,76,77,73,74,51,43,65,30,72,54,92,33,37,75,88,53,84,23,38,86,56,71,68,55,82,62,98,74,81,76,75,23,73,3,45,51,2,92,91,32,44,86,85,5,67,41,36,21,83,52,96,93,84,75,74,94,61,53,72,85,31,87,71,56,80,54,35,64,43,13,5,63,97,82,76,83,3,81,62,33,92,11,93,86,64,37,21,62,30,85,72,34,84,75,18,48,53,95,73,58,44,56,46,59,71,82,19,55,65,63,80,74,33,57,73,78,24,94,72,51,8,55,39,76,64,83,68,86,49,80,7,88,85,32,53,84,37,66,98,99,77,7,85,77,78,65,57,70,84,96,46,13,86,66,75,43,97,89,36,44,59,58,41,74,54,56,55,42,29,92,49,94,88,48,87,43,57,76,53,30,67,58,78,37,66,97,36,32,68,75,47,29,46,49,99,86,56,65,98,50,74,57,77,95,86,68,88,69,81,54,97,76,98,90,42,87,79,75,38,96,25,47,26,67,99,52,80,72,50,58,65,78,5,39,89,80,98,70,47,100,99,67,96,63,88,3,60,86,69,77,76,45,46,56,68,49,48,90,66,61,73,70,59,57,50,51,100,60,89,79,30,98,27,23,78,49,24,5,90,97,74,77,76,88,6,14,19,48,67,69,40,53,71,59,93,91,45,96,87,46,64,73,82,72,83,99,63,33,61,66,4,84,57,21,41,77,92,51,95,62,3,81,62,83,32,100,45,39,91,96,48,57,52,73,84,63,94,78,85,42,36,93,95,47,28,43,72,68,11,89,4,53,88,72,93,52,62,77,84,74,54,22,87,91,32,82,85,67,94,51,63,56,66,92,71,24,28,69,75,86,97,81,65,43,57,74,68,94,92,64,86,72,85,54,61,75,53,33,66,93,91,39,40,73,82,83,97,95,9,63,30,79,74,97,75,95,70,45,63,65,68,3,96,28,66,76,53,55,86,56,42,83,57,71,81,27,88,18,49,25,84,87,97,36,66,85,49,76,39,35,99,94,93,74,43,89,55,18,96,59,16,71,77,95,68,51,52,82,88,23,65,89,95,64,44,57,45,93,84,97,53,77,72,16,60,58,78,86,85,96,68,88,90,79,73,47,67,51,99,81,56,14,10,82,69,87,59,73,98,86,90,47,77,58,89,79,97,48,39,78,28,95,38,63,83,99,65,100,85,75,23,88,67,79,87,30,86,97,90,37,99,64,25,39,80,98,69,96,50,52,58,100,73,43,63,76,91,49,75,94,22,89,100,17,70,85,28,88,67,97,79,40,49,80,48,2,60,87,98,30,5,39,99,77,72,93,62,78,82,95,58,76,92,81,52,62,23,83,42,41,93,82,72,32,21,35,4,61,51,71,37,43,94,63,88,74,49,44,85,7,73,81,14,75,91,93,82,73,53,71,57,52,74,62,87,41,83,72,94,28,32,84,43,86,95,2,44,96,88,51,64,92,34,95,75,63,24,65,85,72,94,82,51,98,49,48,96,84,73,91,81,83,26,71,25,27,11,79,74,23,42,84,67,57,44,95,46,92,63,22,1,7,93,62,85,87,8,73,96,75,97,81,83,82,14,76,65,54,66,48,99,76,85,66,72,65,55,22,92,96,88,49,83,69,47,46,81,44,86,75,50,17,90,87,97,19,51,34,18,93,15,95,77,86,74,76,93,35,84,83,46,92,63,62,67,85,90,33,97,66,94,98,81,75,50,18,89,54,87,36,68,24,47,94,96,95,86,53,99,17,77,83,73,98,100,55,71,76,85,88,65,70,87,56,6,57,49,93,20,90,89,94,97,69,88,14,86,77,91,68,99,100,64,58,59,85,87,78,55,96,79,10,84,23,80,38,60,90,95,89,92,94,89,100,90,98,69,96,95,56,85,59,50,79,58,72,27,49,30,19,40,74,93,68,87,54,63,97,38,64,73,84,80,66,99,90,68,98,88,48,86,59,97,93,79,96,11,27,74,85,53,19,92,89,95,76,70,41,87,77,67);
--       constant post_indx: index_array:=     (44,11,3,4,21,2,22,19,42,14,31,12,35,23,34,15,13,5,41,32,26,52,51,38,29,24,47,33,64,54,33,3,24,3,25,34,12,23,15,5,21,32,10,7,54,22,4,11,6,14,61,42,81,66,28,43,13,52,92,64,14,13,4,5,6,4,22,31,55,4,29,15,63,7,23,12,41,33,43,9,24,11,36,42,62,53,25,44,71,34,28,52,6,14,5,23,7,24,15,5,5,13,11,33,16,26,31,20,22,25,8,54,5,45,18,9,12,41,27,51,6,25,6,14,23,15,17,26,8,16,6,38,7,37,33,59,32,20,13,11,18,6,45,35,19,31,9,27,6,47,7,7,16,7,7,30,59,26,46,8,35,37,17,7,25,15,9,36,13,23,18,24,29,33,34,44,39,12,87,62,8,8,17,16,37,9,28,30,47,25,39,8,18,67,26,27,60,14,75,32,29,24,77,59,20,8,58,8,10,63,18,55,15,37,9,9,19,9,17,40,49,28,39,9,48,9,38,68,29,21,46,9,69,9,20,26,58,10,9,30,28,10,10,19,37,20,10,40,18,39,10,27,50,25,29,26,58,16,10,38,70,49,17,69,54,30,10,87,89,59,29,18,11,20,30,11,17,11,100,38,11,79,19,70,39,58,25,40,35,59,45,66,49,50,11,28,27,60,11,78,12,52,22,14,56,21,94,12,12,15,12,44,32,64,25,55,24,43,31,63,13,81,27,41,61,12,72,83,42,51,14,13,21,13,22,23,13,33,13,13,24,46,16,42,13,26,25,32,13,43,31,52,66,72,63,53,65,54,13,15,14,14,14,23,22,21,73,33,36,16,14,14,14,45,14,17,24,67,20,15,37,14,25,14,51,52,31,63,62,27,15,15,15,24,26,16,15,63,57,15,17,34,66,15,15,15,33,21,23,15,25,27,22,43,41,37,55,73,15,20,16,16,25,28,16,16,16,62,26,36,16,35,37,23,22,45,24,16,38,52,20,39,17,55,42,30,77,47,16,16,19,17,27,17,17,36,17,17,17,17,20,26,25,28,17,56,46,38,34,39,17,17,17,66,47,35,17,57,37,18,27,26,21,18,87,18,25,38,18,18,28,29,45,18,19,18,37,18,44,32,18,18,18,24,47,49,20,39,18,67,28,19,19,37,29,19,22,59,25,38,19,27,55,31,19,69,19,46,19,20,19,36,74,19,26,70,30,48,68,64,30,20,20,39,41,20,20,50,20,20,48,47,29,32,20,20,49,27,20,25,28,20,20,37,38,59,40,65,22,24,21,21,23,29,38,30,50,45,21,21,40,21,28,24,49,21,68,59,33,21,39,66,63,21,60,27,48,21,58,21,22,31,82,22,32,22,25,22,23,33,22,45,22,57,41,22,24,42,43,22,22,56,22,61,22,22,22,64,34,27,46,23,23,31,23,32,24,41,23,52,23,23,23,23,23,23,33,25,23,23,42,55,43,26,62,23,54,53,82,51,34,24,24,24,24,62,24,33,24,24,24,73,25,32,92,31,43,44,24,41,81,26,46,54,24,53,24,24,71,55,25,25,25,25,25,25,34,59,25,33,25,45,32,44,27,25,36,26,64,37,25,30,35,97,25,25,28,74,55,51,27,26,35,26,26,34,26,45,26,31,46,37,26,26,47,26,30,26,28,26,26,26,51,26,38,76,44,77,61,29,27,74,27,27,55,45,28,36,27,46,37,27,32,27,27,47,73,27,34,33,29,27,35,27,27,66,27,58,27,27,28,49,77,28,57,28,76,28,28,28,39,37,70,38,47,61,28,28,28,56,28,58,30,48,55,28,29,28,28,28,38,29,29,29,29,50,58,29,29,55,29,39,79,29,29,30,29,48,29,49,29,60,69,59,37,29,29,47,29,40,30,59,48,47,30,30,39,30,30,30,40,30,30,49,30,30,57,30,37,96,30,65,38,30,30,30,30,60,95,30,31,39,31,40,31,38,45,79,31,31,60,31,57,31,50,49,88,31,70,31,48,59,31,31,31,31,31,90,37,68,32,52,32,41,32,33,32,42,32,81,32,32,32,32,54,61,43,32,51,92,94,35,34,32,46,55,32,64,63,44,42,52,72,33,33,33,62,43,33,41,51,63,33,33,35,33,34,33,44,33,33,64,91,45,82,53,39,54,33,33,34,73,35,43,34,34,34,34,41,42,61,64,34,63,34,34,34,45,39,44,34,54,36,34,57,84,53,46,34,34,35,64,35,35,35,35,46,69,36,44,35,35,35,55,35,45,35,35,52,35,35,35,54,56,79,37,41,35,73,35,37,36,36,36,65,36,88,36,49,36,36,44,36,36,36,45,36,75,40,74,55,36,50,36,36,47,36,46,85,36,37,37,37,37,37,37,37,37,37,48,45,37,37,46,39,37,72,37,38,80,47,37,56,37,37,98,42,37,37,67,38,47,57,38,38,59,67,78,39,38,58,38,38,38,38,38,97,38,75,38,48,54,38,38,85,79,66,38,46,38,39,49,48,56,39,39,39,39,58,40,39,39,46,39,39,39,39,39,55,99,68,59,39,39,66,39,47,39,75,86,40,50,40,49,59,47,40,40,40,40,40,58,40,69,48,40,40,40,68,67,40,57,40,40,60,40,40,40,40,77,41,41,41,59,49,60,41,41,41,41,70,41,48,80,50,41,41,41,41,41,96,93,41,41,79,73,78,41,47,68,42,51,53,45,43,42,62,61,82,42,81,42,42,42,42,52,42,44,83,42,42,48,42,42,71,42,96,63,54,42,45,43,43,72,52,43,62,43,55,51,53,43,61,43,43,43,92,43,73,50,85,43,43,43,83,95,58,43,77,44,63,44,53,44,44,44,44,51,44,54,44,45,83,44,55,47,44,52,44,44,44,44,44,88,44,44,44,46,74,58,45,64,45,45,46,54,45,45,45,45,45,93,49,45,45,45,53,45,69,50,84,52,45,45,65,74,57,81,45,45,55,46,48,46,46,85,72,54,46,46,46,53,46,66,46,97,46,46,95,46,56,52,84,46,46,46,65,46,76,46,47,47,54,47,55,47,53,47,56,47,96,47,47,47,82,92,47,67,47,57,48,47,47,49,63,47,66,78,84,87,48,48,48,57,48,48,48,48,48,48,48,67,60,48,74,48,48,48,58,77,49,50,84,48,85,66,78,68,54,89,49,49,68,78,49,79,50,49,49,49,49,49,49,52,49,49,49,49,49,66,49,49,58,69,57,98,49,72,60,90,50,50,50,69,59,50,50,50,50,50,50,50,79,50,76,57,50,50,50,53,50,58,50,50,50,86,50,97,50,65,51,79,80,67,51,60,51,59,78,51,69,51,51,51,51,58,51,57,51,51,51,51,70,51,51,51,51,51,55,51,53,62,84,52,71,52,52,52,52,74,52,52,61,81,63,52,92,52,55,54,52,83,52,72,75,52,52,95,76,64,62,53,61,85,55,72,53,78,53,82,53,81,80,53,64,53,53,71,77,74,54,73,53,92,57,84,53,63,53,53,56,63,54,54,54,54,65,54,85,54,54,54,73,54,54,81,62,54,91,54,83,54,72,54,64,61,54,57,92,54,55,56,91,55,64,65,55,84,74,55,55,81,75,55,55,55,70,55,93,57,63,85,55,55,55,61,55,55,55,55,65,56,57,56,56,56,64,56,71,56,83,63,56,56,56,56,73,75,85,56,56,66,56,68,56,56,56,56,56,56,57,57,66,57,58,86,57,78,89,57,57,60,57,57,57,57,57,77,57,57,57,69,57,76,57,59,57,98,57,74,58,68,67,58,70,69,59,64,77,58,58,86,83,58,76,58,58,60,80,66,75,61,63,58,88,58,58,58,98,78,68,59,59,59,67,59,59,59,59,59,59,60,80,59,88,97,78,70,59,87,59,74,64,77,59,59,69,59,59,86,60,79,60,60,60,69,89,94,96,60,60,60,60,68,90,100,60,60,60,60,60,88,99,80,60,60,65,70,98,66,61,67,61,61,61,90,61,80,100,70,96,79,61,75,61,61,69,68,61,61,61,61,76,78,88,61,77,61,61,61,62,63,62,71,81,73,62,62,62,83,72,75,91,82,62,64,62,62,62,65,92,66,62,87,62,62,95,62,62,62,64,63,73,63,72,63,82,63,63,63,63,63,92,74,63,65,81,63,63,63,71,95,63,63,63,96,63,63,63,63,64,64,93,73,64,64,66,64,64,71,64,65,64,84,64,75,64,74,64,96,83,72,64,64,64,64,64,64,64,64,65,65,71,75,65,65,65,66,65,85,96,65,65,84,83,74,87,73,94,65,76,65,65,65,77,65,65,65,65,65,76,95,66,66,83,96,75,66,66,66,66,66,69,73,70,66,78,66,67,86,66,66,66,66,66,66,66,85,66,66,67,67,86,67,67,76,67,67,68,67,75,67,67,85,67,67,67,77,98,67,69,67,67,71,79,97,67,99,67,67,68,68,77,68,68,87,68,68,68,97,68,68,68,89,68,68,68,76,100,68,68,84,68,79,96,68,68,68,68,69,69,69,69,89,69,98,69,69,78,76,69,69,69,69,69,69,69,69,77,69,69,69,69,79,69,70,69,87,88,69,79,89,70,70,70,99,70,70,98,70,70,80,70,86,90,78,70,70,70,70,70,73,70,70,70,70,70,97,70,70,100,71,89,71,71,79,71,71,71,71,71,99,71,80,71,90,86,71,71,71,71,98,71,71,71,87,71,71,84,77,72,91,72,72,72,72,72,72,72,81,72,85,82,76,72,72,83,73,74,72,72,72,72,93,72,92,72,72,72,72,92,73,94,73,75,82,73,81,73,73,73,83,73,73,73,73,73,73,73,73,95,73,73,73,73,73,93,73,73,73,74,74,74,94,74,74,74,74,74,74,76,82,86,84,74,74,93,74,74,85,74,83,81,75,74,74,74,74,74,92,75,75,75,75,75,76,75,75,94,75,83,77,90,75,80,75,84,75,85,91,75,75,75,75,75,75,81,75,88,75,85,82,78,97,76,95,77,76,81,76,76,76,76,76,84,76,76,76,79,76,76,76,76,96,87,76,76,76,86,76,77,77,77,87,96,86,77,93,83,77,77,77,94,88,77,77,77,77,77,95,77,77,77,77,77,77,77,97,98,84,78,89,78,95,78,78,78,78,96,78,87,88,78,78,97,78,78,78,79,78,78,78,78,78,80,86,78,94,78,90,79,87,86,99,88,79,89,80,79,79,79,79,79,79,98,97,79,79,79,100,96,79,79,79,79,79,90,79,79,79,89,80,80,80,80,99,90,80,80,80,80,80,80,80,80,85,80,100,80,80,80,87,98,97,94,80,80,86,80,80,81,81,81,89,84,90,81,81,81,99,81,100,98,81,81,81,81,81,81,81,81,81,97,81,81,87,81,81,81,81,82,82,91,92,82,82,82,82,93,90,86,82,82,96,82,82,85,83,82,82,82,82,84,82,94,82,82,82,82,88,92,83,83,83,91,83,94,83,83,87,83,83,93,83,83,83,83,85,83,83,83,84,86,90,83,83,83,83,83,83,84,84,85,84,84,93,94,84,84,84,84,84,84,88,92,96,84,84,91,84,84,84,84,84,84,95,84,97,100,84,85,85,86,85,85,85,93,92,85,85,88,95,85,85,97,94,85,85,85,85,85,85,85,85,85,85,85,85,85,85,86,86,87,86,86,95,94,86,86,86,86,90,86,86,86,86,86,96,86,86,86,86,97,86,86,99,86,86,86,86,87,87,87,96,87,98,87,87,87,87,87,95,87,87,87,97,87,87,92,87,87,87,87,87,87,88,87,87,87,87,88,88,88,88,88,88,88,97,88,98,88,88,89,94,88,88,88,88,96,88,88,88,100,88,88,88,99,92,88,88,96,89,89,89,89,89,89,95,89,89,90,89,89,98,89,89,99,89,89,97,89,100,89,89,89,89,89,89,89,89,90,90,90,98,99,90,90,90,90,100,90,90,90,90,90,90,90,90,90,90,97,90,90,90,93,96,90,90,90,90,91,91,91,91,91,91,91,91,91,100,91,91,91,91,91,91,91,96,91,91,98,91,97,99,91,91,91,91,91,91,92,92,92,92,92,92,92,92,92,97,92,96,92,93,99,92,92,94,92,92,92,92,95,92,92,92,92,92,92,92,95,93,94,93,93,93,93,93,93,93,93,96,93,93,97,93,93,93,93,93,93,93,93,93,93,93,100,93,93,93,94,94,94,94,94,96,94,94,94,94,95,94,94,97,94,94,94,94,94,98,94,94,94,94,94,94,94,94,94,94,95,95,95,95,95,95,95,95,95,95,95,97,95,95,95,95,95,95,95,95,100,95,95,95,95,95,96,95,95,99,97,96,96,96,96,96,96,96,96,96,96,96,96,100,96,96,96,96,96,96,98,96,96,96,96,96,96,96,96,96,97,97,97,97,97,97,97,97,98,97,97,97,97,97,97,97,97,97,97,97,99,97,97,97,97,97,97,97,97,97,98,98,98,98,98,98,98,98,98,98,98,98,98,98,99,98,98,98,98,98,98,100,98,98,98,98,98,98,98,98,99,99,99,99,99,99,99,99,100,99,99,99,99,99,99,99,99,99,99,99,99,99,99,99,99,99,99,99,99,99,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100,100);
constant post_indx: index_array:=(21 ,
4  ,
33 ,
11 ,
2  ,
12 ,
13 ,
22 ,
25 ,
23 ,
3  ,
32 ,
14 ,
6  ,
42 ,
5  ,
41 ,
51 ,
31 ,
8  ,
12 ,
13 ,
3  ,
21 ,
1  ,
5  ,
27 ,
14 ,
4  ,
22 ,
11 ,
54 ,
41 ,
23 ,
33 ,
28 ,
32 ,
24 ,
6  ,
43 ,
5  ,
2  ,
13 ,
4  ,
23 ,
12 ,
24 ,
25 ,
1  ,
15 ,
35 ,
6  ,
53 ,
52 ,
22 ,
14 ,
16 ,
11 ,
33 ,
21 ,
5  ,
3  ,
16 ,
14 ,
25 ,
15 ,
26 ,
17 ,
23 ,
2  ,
34 ,
11 ,
22 ,
6  ,
24 ,
12 ,
1  ,
7  ,
13 ,
32 ,
23 ,
4  ,
26 ,
16 ,
35 ,
15 ,
3  ,
6  ,
8  ,
25 ,
7  ,
13 ,
14 ,
24 ,
36 ,
2  ,
17 ,
27 ,
57 ,
45 ,
5  ,
7  ,
34 ,
16 ,
10 ,
26 ,
14 ,
17 ,
18 ,
42 ,
4  ,
28 ,
15 ,
29 ,
8  ,
23 ,
36 ,
30 ,
56 ,
3  ,
17 ,
5  ,
8  ,
19 ,
6  ,
47 ,
30 ,
28 ,
9  ,
45 ,
14 ,
3  ,
18 ,
38 ,
16 ,
37 ,
25 ,
26 ,
27 ,
60 ,
18 ,
27 ,
10 ,
9  ,
6  ,
36 ,
20 ,
7  ,
16 ,
28 ,
40 ,
17 ,
19 ,
47 ,
39 ,
44 ,
37 ,
5  ,
26 ,
38 ,
8  ,
19 ,
10 ,
39 ,
29 ,
20 ,
38 ,
18 ,
17 ,
7  ,
15 ,
30 ,
16 ,
49 ,
27 ,
6  ,
28 ,
78 ,
35 ,
37 ,
29 ,
9  ,
20 ,
30 ,
19 ,
17 ,
18 ,
8  ,
40 ,
16 ,
28 ,
7  ,
47 ,
39 ,
59 ,
27 ,
6  ,
50 ,
67 ,
26 ,
12 ,
23 ,
1  ,
21 ,
13 ,
31 ,
2  ,
22 ,
42 ,
41 ,
4  ,
62 ,
61 ,
15 ,
33 ,
43 ,
14 ,
3  ,
29 ,
32 ,
32 ,
43 ,
13 ,
22 ,
2  ,
1  ,
3  ,
25 ,
14 ,
23 ,
24 ,
11 ,
4  ,
31 ,
21 ,
42 ,
33 ,
15 ,
16 ,
65 ,
23 ,
14 ,
24 ,
4  ,
33 ,
3  ,
12 ,
25 ,
34 ,
22 ,
44 ,
1  ,
21 ,
11 ,
43 ,
32 ,
16 ,
15 ,
56 ,
2  ,
3  ,
21 ,
13 ,
12 ,
15 ,
4  ,
24 ,
22 ,
31 ,
34 ,
5  ,
33 ,
23 ,
25 ,
1  ,
11 ,
35 ,
62 ,
6  ,
43 ,
14 ,
25 ,
17 ,
5  ,
24 ,
13 ,
35 ,
4  ,
36 ,
48 ,
16 ,
45 ,
26 ,
6  ,
3  ,
27 ,
44 ,
33 ,
22 ,
46 ,
6  ,
15 ,
14 ,
24 ,
36 ,
18 ,
5  ,
17 ,
19 ,
25 ,
8  ,
27 ,
10 ,
37 ,
20 ,
26 ,
35 ,
7  ,
57 ,
45 ,
26 ,
15 ,
20 ,
16 ,
27 ,
19 ,
37 ,
7  ,
6  ,
25 ,
18 ,
14 ,
36 ,
8  ,
9  ,
5  ,
38 ,
29 ,
28 ,
45 ,
48 ,
27 ,
17 ,
8  ,
19 ,
10 ,
29 ,
9  ,
28 ,
26 ,
6  ,
37 ,
15 ,
59 ,
35 ,
16 ,
36 ,
5  ,
7  ,
38 ,
30 ,
18 ,
39 ,
20 ,
29 ,
28 ,
40 ,
16 ,
37 ,
8  ,
9  ,
7  ,
5  ,
10 ,
17 ,
49 ,
36 ,
38 ,
27 ,
88 ,
29 ,
30 ,
40 ,
50 ,
38 ,
19 ,
17 ,
10 ,
48 ,
18 ,
28 ,
27 ,
9  ,
8  ,
7  ,
60 ,
59 ,
37 ,
49 ,
39 ,
22 ,
31 ,
11 ,
53 ,
32 ,
23 ,
41 ,
12 ,
13 ,
42 ,
1  ,
44 ,
2  ,
33 ,
43 ,
3  ,
51 ,
14 ,
52 ,
24 ,
21 ,
33 ,
31 ,
12 ,
23 ,
2  ,
52 ,
3  ,
25 ,
11 ,
13 ,
34 ,
32 ,
1  ,
4  ,
42 ,
53 ,
24 ,
26 ,
44 ,
58 ,
24 ,
33 ,
32 ,
22 ,
28 ,
5  ,
21 ,
13 ,
53 ,
83 ,
43 ,
14 ,
4  ,
26 ,
36 ,
25 ,
61 ,
34 ,
12 ,
61 ,
34 ,
23 ,
14 ,
25 ,
31 ,
26 ,
22 ,
42 ,
41 ,
27 ,
35 ,
56 ,
75 ,
15 ,
87 ,
33 ,
12 ,
4  ,
7  ,
15 ,
35 ,
53 ,
14 ,
45 ,
22 ,
16 ,
4  ,
36 ,
34 ,
5  ,
27 ,
24 ,
26 ,
46 ,
38 ,
43 ,
12 ,
23 ,
55 ,
24 ,
25 ,
36 ,
47 ,
17 ,
46 ,
16 ,
28 ,
34 ,
27 ,
37 ,
15 ,
35 ,
5  ,
18 ,
43 ,
76 ,
45 ,
32 ,
48 ,
26 ,
47 ,
57 ,
37 ,
58 ,
25 ,
28 ,
36 ,
16 ,
17 ,
18 ,
29 ,
5  ,
45 ,
35 ,
6  ,
46 ,
38 ,
40 ,
19 ,
27 ,
18 ,
38 ,
8  ,
48 ,
29 ,
26 ,
19 ,
39 ,
9  ,
30 ,
6  ,
14 ,
49 ,
45 ,
68 ,
70 ,
58 ,
40 ,
17 ,
39 ,
24 ,
19 ,
30 ,
20 ,
10 ,
28 ,
68 ,
26 ,
58 ,
27 ,
38 ,
50 ,
49 ,
37 ,
60 ,
35 ,
59 ,
40 ,
9  ,
29 ,
40 ,
20 ,
28 ,
50 ,
60 ,
59 ,
38 ,
39 ,
10 ,
18 ,
27 ,
9  ,
68 ,
80 ,
19 ,
26 ,
17 ,
47 ,
48 ,
22 ,
51 ,
42 ,
11 ,
21 ,
41 ,
61 ,
33 ,
53 ,
32 ,
23 ,
34 ,
83 ,
2  ,
1  ,
12 ,
43 ,
62 ,
63 ,
35 ,
34 ,
31 ,
42 ,
22 ,
43 ,
5  ,
41 ,
21 ,
64 ,
44 ,
52 ,
33 ,
63 ,
14 ,
51 ,
12 ,
13 ,
23 ,
36 ,
15 ,
43 ,
32 ,
13 ,
34 ,
52 ,
23 ,
22 ,
31 ,
53 ,
35 ,
71 ,
24 ,
46 ,
20 ,
44 ,
42 ,
25 ,
45 ,
64 ,
21 ,
35 ,
33 ,
38 ,
54 ,
24 ,
53 ,
44 ,
31 ,
14 ,
74 ,
56 ,
23 ,
37 ,
27 ,
45 ,
25 ,
62 ,
43 ,
42 ,
65 ,
25 ,
45 ,
57 ,
36 ,
24 ,
38 ,
56 ,
34 ,
22 ,
28 ,
47 ,
37 ,
55 ,
31 ,
21 ,
33 ,
41 ,
14 ,
76 ,
48 ,
26 ,
46 ,
37 ,
38 ,
35 ,
15 ,
16 ,
27 ,
56 ,
34 ,
25 ,
47 ,
39 ,
24 ,
32 ,
33 ,
7  ,
43 ,
23 ,
6  ,
36 ,
27 ,
47 ,
56 ,
26 ,
38 ,
46 ,
15 ,
39 ,
17 ,
77 ,
35 ,
58 ,
48 ,
28 ,
57 ,
18 ,
34 ,
23 ,
45 ,
68 ,
59 ,
49 ,
8  ,
37 ,
40 ,
28 ,
29 ,
27 ,
18 ,
48 ,
36 ,
39 ,
70 ,
17 ,
7  ,
6  ,
47 ,
25 ,
78 ,
48 ,
29 ,
49 ,
50 ,
40 ,
38 ,
28 ,
57 ,
16 ,
9  ,
58 ,
59 ,
27 ,
37 ,
19 ,
26 ,
80 ,
30 ,
60 ,
20 ,
50 ,
20 ,
39 ,
30 ,
38 ,
19 ,
29 ,
90 ,
26 ,
49 ,
60 ,
76 ,
70 ,
48 ,
10 ,
28 ,
57 ,
47 ,
59 ,
89 ,
42 ,
43 ,
31 ,
33 ,
62 ,
51 ,
22 ,
32 ,
61 ,
52 ,
21 ,
71 ,
53 ,
11 ,
63 ,
73 ,
2  ,
44 ,
16 ,
45 ,
52 ,
41 ,
53 ,
63 ,
43 ,
62 ,
32 ,
44 ,
21 ,
31 ,
51 ,
61 ,
22 ,
33 ,
81 ,
71 ,
72 ,
55 ,
12 ,
83 ,
33 ,
53 ,
42 ,
3  ,
34 ,
13 ,
14 ,
32 ,
64 ,
41 ,
62 ,
44 ,
31 ,
85 ,
73 ,
12 ,
22 ,
24 ,
63 ,
54 ,
34 ,
83 ,
24 ,
42 ,
54 ,
66 ,
41 ,
43 ,
56 ,
55 ,
68 ,
84 ,
64 ,
45 ,
46 ,
33 ,
53 ,
12 ,
74 ,
63 ,
55 ,
95 ,
23 ,
78 ,
35 ,
44 ,
65 ,
43 ,
42 ,
46 ,
63 ,
25 ,
56 ,
48 ,
36 ,
47 ,
85 ,
33 ,
57 ,
54 ,
37 ,
89 ,
45 ,
56 ,
38 ,
47 ,
66 ,
36 ,
26 ,
35 ,
69 ,
24 ,
48 ,
67 ,
44 ,
55 ,
43 ,
17 ,
77 ,
49 ,
77 ,
27 ,
56 ,
49 ,
68 ,
39 ,
55 ,
57 ,
16 ,
44 ,
17 ,
37 ,
48 ,
65 ,
59 ,
36 ,
46 ,
45 ,
7  ,
67 ,
39 ,
49 ,
58 ,
47 ,
60 ,
28 ,
68 ,
38 ,
27 ,
59 ,
50 ,
37 ,
78 ,
26 ,
40 ,
55 ,
66 ,
69 ,
57 ,
67 ,
50 ,
70 ,
39 ,
38 ,
58 ,
59 ,
36 ,
48 ,
57 ,
69 ,
30 ,
78 ,
29 ,
99 ,
47 ,
18 ,
46 ,
19 ,
67 ,
68 ,
49 ,
30 ,
40 ,
87 ,
65 ,
60 ,
48 ,
59 ,
78 ,
70 ,
39 ,
47 ,
57 ,
46 ,
36 ,
19 ,
8  ,
25 ,
69 ,
80 ,
52 ,
61 ,
41 ,
71 ,
81 ,
21 ,
62 ,
42 ,
31 ,
12 ,
63 ,
57 ,
82 ,
83 ,
35 ,
72 ,
43 ,
46 ,
53 ,
54 ,
53 ,
42 ,
62 ,
32 ,
54 ,
61 ,
72 ,
51 ,
41 ,
71 ,
63 ,
64 ,
66 ,
55 ,
34 ,
31 ,
73 ,
46 ,
65 ,
81 ,
52 ,
55 ,
45 ,
64 ,
73 ,
41 ,
54 ,
63 ,
43 ,
97 ,
72 ,
62 ,
51 ,
81 ,
33 ,
22 ,
23 ,
3  ,
67 ,
12 ,
44 ,
45 ,
64 ,
62 ,
55 ,
67 ,
53 ,
51 ,
52 ,
42 ,
43 ,
12 ,
58 ,
74 ,
76 ,
56 ,
63 ,
68 ,
72 ,
24 ,
57 ,
67 ,
37 ,
53 ,
65 ,
35 ,
22 ,
45 ,
54 ,
56 ,
24 ,
74 ,
75 ,
40 ,
52 ,
47 ,
25 ,
73 ,
43 ,
34 ,
57 ,
27 ,
55 ,
66 ,
65 ,
46 ,
54 ,
58 ,
43 ,
77 ,
16 ,
26 ,
68 ,
87 ,
44 ,
36 ,
47 ,
76 ,
53 ,
86 ,
46 ,
47 ,
56 ,
67 ,
87 ,
66 ,
37 ,
79 ,
58 ,
59 ,
55 ,
86 ,
35 ,
68 ,
65 ,
48 ,
27 ,
26 ,
54 ,
45 ,
57 ,
38 ,
47 ,
60 ,
30 ,
46 ,
59 ,
40 ,
78 ,
56 ,
68 ,
20 ,
85 ,
49 ,
69 ,
28 ,
48 ,
87 ,
17 ,
77 ,
69 ,
57 ,
60 ,
39 ,
49 ,
99 ,
58 ,
80 ,
56 ,
70 ,
98 ,
29 ,
40 ,
68 ,
48 ,
88 ,
55 ,
50 ,
90 ,
28 ,
49 ,
70 ,
79 ,
59 ,
47 ,
68 ,
39 ,
58 ,
50 ,
48 ,
69 ,
56 ,
28 ,
30 ,
80 ,
67 ,
40 ,
66 ,
78 ,
88 ,
51 ,
73 ,
62 ,
71 ,
81 ,
53 ,
52 ,
92 ,
31 ,
41 ,
82 ,
72 ,
63 ,
74 ,
42 ,
91 ,
85 ,
83 ,
23 ,
64 ,
61 ,
72 ,
63 ,
82 ,
64 ,
91 ,
73 ,
52 ,
74 ,
45 ,
25 ,
42 ,
53 ,
32 ,
51 ,
92 ,
71 ,
55 ,
75 ,
43 ,
65 ,
62 ,
72 ,
44 ,
43 ,
74 ,
61 ,
64 ,
83 ,
73 ,
71 ,
53 ,
67 ,
93 ,
57 ,
82 ,
84 ,
95 ,
55 ,
81 ,
63 ,
84 ,
65 ,
53 ,
92 ,
93 ,
74 ,
34 ,
66 ,
54 ,
94 ,
73 ,
43 ,
78 ,
55 ,
67 ,
77 ,
68 ,
51 ,
45 ,
73 ,
64 ,
66 ,
85 ,
55 ,
75 ,
33 ,
67 ,
83 ,
44 ,
86 ,
46 ,
76 ,
45 ,
87 ,
63 ,
57 ,
54 ,
47 ,
53 ,
76 ,
34 ,
67 ,
65 ,
15 ,
77 ,
46 ,
56 ,
59 ,
75 ,
86 ,
55 ,
85 ,
74 ,
64 ,
89 ,
21 ,
72 ,
57 ,
63 ,
77 ,
53 ,
76 ,
97 ,
66 ,
47 ,
46 ,
55 ,
57 ,
69 ,
68 ,
64 ,
27 ,
58 ,
49 ,
65 ,
87 ,
59 ,
78 ,
89 ,
77 ,
67 ,
58 ,
76 ,
60 ,
59 ,
78 ,
57 ,
69 ,
47 ,
88 ,
79 ,
70 ,
97 ,
99 ,
65 ,
74 ,
98 ,
48 ,
66 ,
68 ,
80 ,
70 ,
59 ,
79 ,
89 ,
50 ,
60 ,
67 ,
48 ,
78 ,
49 ,
65 ,
37 ,
57 ,
38 ,
58 ,
56 ,
98 ,
20 ,
49 ,
66 ,
60 ,
100,
69 ,
59 ,
85 ,
80 ,
77 ,
50 ,
20 ,
78 ,
79 ,
90 ,
67 ,
30 ,
68 ,
88 ,
99 ,
58 ,
72 ,
81 ,
85 ,
74 ,
82 ,
73 ,
91 ,
62 ,
42 ,
63 ,
61 ,
67 ,
51 ,
43 ,
92 ,
83 ,
41 ,
52 ,
93 ,
31 ,
62 ,
71 ,
52 ,
24 ,
73 ,
81 ,
82 ,
61 ,
47 ,
63 ,
51 ,
42 ,
83 ,
75 ,
45 ,
53 ,
91 ,
33 ,
46 ,
74 ,
72 ,
63 ,
74 ,
54 ,
52 ,
93 ,
83 ,
75 ,
62 ,
85 ,
82 ,
64 ,
71 ,
44 ,
56 ,
84 ,
43 ,
81 ,
53 ,
94 ,
84 ,
65 ,
54 ,
73 ,
76 ,
75 ,
94 ,
85 ,
72 ,
48 ,
83 ,
62 ,
64 ,
63 ,
77 ,
98 ,
34 ,
71 ,
82 ,
44 ,
65 ,
55 ,
85 ,
86 ,
74 ,
44 ,
96 ,
73 ,
84 ,
95 ,
77 ,
76 ,
94 ,
62 ,
97 ,
66 ,
99 ,
54 ,
57 ,
56 ,
66 ,
78 ,
75 ,
87 ,
99 ,
86 ,
77 ,
39 ,
74 ,
54 ,
95 ,
85 ,
47 ,
35 ,
23 ,
64 ,
55 ,
82 ,
56 ,
80 ,
76 ,
78 ,
69 ,
67 ,
66 ,
59 ,
95 ,
68 ,
35 ,
74 ,
88 ,
97 ,
58 ,
57 ,
27 ,
98 ,
79 ,
87 ,
96 ,
80 ,
58 ,
79 ,
77 ,
88 ,
74 ,
76 ,
48 ,
90 ,
80 ,
14 ,
98 ,
68 ,
69 ,
67 ,
87 ,
97 ,
35 ,
70 ,
89 ,
66 ,
97 ,
68 ,
78 ,
99 ,
80 ,
100,
98 ,
60 ,
67 ,
76 ,
89 ,
69 ,
59 ,
70 ,
30 ,
77 ,
88 ,
75 ,
49 ,
58 ,
60 ,
100,
79 ,
70 ,
68 ,
89 ,
88 ,
48 ,
90 ,
77 ,
69 ,
78 ,
76 ,
75 ,
86 ,
59 ,
27 ,
98 ,
12 ,
20 ,
71 ,
91 ,
92 ,
82 ,
93 ,
61 ,
63 ,
51 ,
53 ,
42 ,
73 ,
52 ,
83 ,
43 ,
72 ,
84 ,
74 ,
96 ,
44 ,
54 ,
92 ,
85 ,
72 ,
83 ,
62 ,
52 ,
81 ,
34 ,
94 ,
84 ,
93 ,
73 ,
91 ,
74 ,
63 ,
71 ,
61 ,
86 ,
53 ,
42 ,
84 ,
53 ,
74 ,
94 ,
82 ,
93 ,
72 ,
92 ,
63 ,
52 ,
85 ,
73 ,
87 ,
65 ,
81 ,
61 ,
43 ,
62 ,
95 ,
98 ,
82 ,
83 ,
64 ,
93 ,
75 ,
74 ,
94 ,
85 ,
96 ,
95 ,
86 ,
54 ,
65 ,
73 ,
76 ,
62 ,
55 ,
72 ,
67 ,
63 ,
96 ,
84 ,
92 ,
63 ,
56 ,
95 ,
86 ,
55 ,
76 ,
74 ,
88 ,
83 ,
75 ,
94 ,
77 ,
67 ,
62 ,
65 ,
64 ,
97 ,
96 ,
76 ,
87 ,
66 ,
88 ,
95 ,
85 ,
97 ,
77 ,
68 ,
90 ,
57 ,
75 ,
28 ,
74 ,
84 ,
98 ,
45 ,
93 ,
56 ,
88 ,
91 ,
77 ,
96 ,
76 ,
86 ,
68 ,
89 ,
85 ,
97 ,
98 ,
99 ,
79 ,
67 ,
69 ,
90 ,
75 ,
47 ,
78 ,
84 ,
90 ,
98 ,
78 ,
87 ,
68 ,
99 ,
86 ,
94 ,
66 ,
59 ,
89 ,
69 ,
100,
85 ,
97 ,
67 ,
70 ,
84 ,
65 ,
80 ,
79 ,
90 ,
87 ,
88 ,
99 ,
97 ,
100,
78 ,
69 ,
59 ,
76 ,
68 ,
80 ,
77 ,
58 ,
66 ,
98 ,
67 ,
96 ,
86 ,
79 ,
100,
89 ,
80 ,
88 ,
76 ,
87 ,
99 ,
66 ,
68 ,
58 ,
70 ,
69 ,
78 ,
86 ,
60 ,
59 ,
98 ,
77 ,
97 ,
82 ,
71 ,
92 ,
81 ,
64 ,
93 ,
84 ,
72 ,
94 ,
83 ,
63 ,
73 ,
62 ,
96 ,
61 ,
95 ,
52 ,
74 ,
51 ,
53 ,
93 ,
91 ,
82 ,
83 ,
84 ,
55 ,
94 ,
71 ,
95 ,
86 ,
52 ,
44 ,
73 ,
64 ,
72 ,
81 ,
63 ,
61 ,
62 ,
85 ,
81 ,
82 ,
92 ,
83 ,
97 ,
94 ,
73 ,
65 ,
91 ,
72 ,
84 ,
85 ,
95 ,
75 ,
98 ,
53 ,
88 ,
74 ,
96 ,
63 ,
73 ,
84 ,
74 ,
93 ,
95 ,
96 ,
75 ,
85 ,
62 ,
97 ,
92 ,
72 ,
81 ,
83 ,
64 ,
99 ,
82 ,
54 ,
91 ,
87 ,
85 ,
96 ,
84 ,
92 ,
88 ,
94 ,
86 ,
97 ,
75 ,
77 ,
81 ,
93 ,
99 ,
74 ,
65 ,
83 ,
71 ,
87 ,
56 ,
55 ,
97 ,
86 ,
94 ,
54 ,
75 ,
95 ,
76 ,
74 ,
98 ,
85 ,
87 ,
65 ,
56 ,
66 ,
78 ,
57 ,
88 ,
37 ,
83 ,
99 ,
88 ,
85 ,
96 ,
98 ,
78 ,
77 ,
95 ,
58 ,
99 ,
87 ,
86 ,
90 ,
92 ,
89 ,
67 ,
94 ,
68 ,
60 ,
76 ,
75 ,
99 ,
87 ,
78 ,
89 ,
100,
96 ,
97 ,
95 ,
86 ,
68 ,
88 ,
80 ,
70 ,
77 ,
79 ,
74 ,
57 ,
90 ,
66 ,
69 ,
89 ,
100,
98 ,
88 ,
68 ,
79 ,
97 ,
87 ,
67 ,
90 ,
69 ,
80 ,
95 ,
78 ,
59 ,
77 ,
96 ,
50 ,
76 ,
85 ,
99 ,
98 ,
90 ,
80 ,
79 ,
89 ,
70 ,
69 ,
76 ,
78 ,
88 ,
59 ,
84 ,
87 ,
97 ,
95 ,
94 ,
77 ,
60 ,
39 );

end package wm_package; 
-- Package Body Section
package body wm_package is
 
  
end package body wm_package;
