

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


package wm_package is

constant  Data_Width: integer:=32;
constant  shift_param:integer:=16;
constant  NN_size:integer:=100;
constant  connection_size:integer:=20;
constant  astro_size:integer:=9;

 type index_array is array (0 to NN_size*connection_size-1) of integer range 0 to 100;------------------ array for saving neuron outputs
 
constant post_indx: index_array:=(21 ,
4  ,
33 ,
11 ,
2  ,
12 ,
13 ,
22 ,
25 ,
23 ,
3  ,
32 ,
14 ,
6  ,
42 ,
5  ,
41 ,
51 ,
31 ,
8  ,
12 ,
13 ,
3  ,
21 ,
1  ,
5  ,
27 ,
14 ,
4  ,
22 ,
11 ,
54 ,
41 ,
23 ,
33 ,
28 ,
32 ,
24 ,
6  ,
43 ,
5  ,
2  ,
13 ,
4  ,
23 ,
12 ,
24 ,
25 ,
1  ,
15 ,
35 ,
6  ,
53 ,
52 ,
22 ,
14 ,
16 ,
11 ,
33 ,
21 ,
5  ,
3  ,
16 ,
14 ,
25 ,
15 ,
26 ,
17 ,
23 ,
2  ,
34 ,
11 ,
22 ,
6  ,
24 ,
12 ,
1  ,
7  ,
13 ,
32 ,
23 ,
4  ,
26 ,
16 ,
35 ,
15 ,
3  ,
6  ,
8  ,
25 ,
7  ,
13 ,
14 ,
24 ,
36 ,
2  ,
17 ,
27 ,
57 ,
45 ,
5  ,
7  ,
34 ,
16 ,
10 ,
26 ,
14 ,
17 ,
18 ,
42 ,
4  ,
28 ,
15 ,
29 ,
8  ,
23 ,
36 ,
30 ,
56 ,
3  ,
17 ,
5  ,
8  ,
19 ,
6  ,
47 ,
30 ,
28 ,
9  ,
45 ,
14 ,
3  ,
18 ,
38 ,
16 ,
37 ,
25 ,
26 ,
27 ,
60 ,
18 ,
27 ,
10 ,
9  ,
6  ,
36 ,
20 ,
7  ,
16 ,
28 ,
40 ,
17 ,
19 ,
47 ,
39 ,
44 ,
37 ,
5  ,
26 ,
38 ,
8  ,
19 ,
10 ,
39 ,
29 ,
20 ,
38 ,
18 ,
17 ,
7  ,
15 ,
30 ,
16 ,
49 ,
27 ,
6  ,
28 ,
78 ,
35 ,
37 ,
29 ,
9  ,
20 ,
30 ,
19 ,
17 ,
18 ,
8  ,
40 ,
16 ,
28 ,
7  ,
47 ,
39 ,
59 ,
27 ,
6  ,
50 ,
67 ,
26 ,
12 ,
23 ,
1  ,
21 ,
13 ,
31 ,
2  ,
22 ,
42 ,
41 ,
4  ,
62 ,
61 ,
15 ,
33 ,
43 ,
14 ,
3  ,
29 ,
32 ,
32 ,
43 ,
13 ,
22 ,
2  ,
1  ,
3  ,
25 ,
14 ,
23 ,
24 ,
11 ,
4  ,
31 ,
21 ,
42 ,
33 ,
15 ,
16 ,
65 ,
23 ,
14 ,
24 ,
4  ,
33 ,
3  ,
12 ,
25 ,
34 ,
22 ,
44 ,
1  ,
21 ,
11 ,
43 ,
32 ,
16 ,
15 ,
56 ,
2  ,
3  ,
21 ,
13 ,
12 ,
15 ,
4  ,
24 ,
22 ,
31 ,
34 ,
5  ,
33 ,
23 ,
25 ,
1  ,
11 ,
35 ,
62 ,
6  ,
43 ,
14 ,
25 ,
17 ,
5  ,
24 ,
13 ,
35 ,
4  ,
36 ,
48 ,
16 ,
45 ,
26 ,
6  ,
3  ,
27 ,
44 ,
33 ,
22 ,
46 ,
6  ,
15 ,
14 ,
24 ,
36 ,
18 ,
5  ,
17 ,
19 ,
25 ,
8  ,
27 ,
10 ,
37 ,
20 ,
26 ,
35 ,
7  ,
57 ,
45 ,
26 ,
15 ,
20 ,
16 ,
27 ,
19 ,
37 ,
7  ,
6  ,
25 ,
18 ,
14 ,
36 ,
8  ,
9  ,
5  ,
38 ,
29 ,
28 ,
45 ,
48 ,
27 ,
17 ,
8  ,
19 ,
10 ,
29 ,
9  ,
28 ,
26 ,
6  ,
37 ,
15 ,
59 ,
35 ,
16 ,
36 ,
5  ,
7  ,
38 ,
30 ,
18 ,
39 ,
20 ,
29 ,
28 ,
40 ,
16 ,
37 ,
8  ,
9  ,
7  ,
5  ,
10 ,
17 ,
49 ,
36 ,
38 ,
27 ,
88 ,
29 ,
30 ,
40 ,
50 ,
38 ,
19 ,
17 ,
10 ,
48 ,
18 ,
28 ,
27 ,
9  ,
8  ,
7  ,
60 ,
59 ,
37 ,
49 ,
39 ,
22 ,
31 ,
11 ,
53 ,
32 ,
23 ,
41 ,
12 ,
13 ,
42 ,
1  ,
44 ,
2  ,
33 ,
43 ,
3  ,
51 ,
14 ,
52 ,
24 ,
21 ,
33 ,
31 ,
12 ,
23 ,
2  ,
52 ,
3  ,
25 ,
11 ,
13 ,
34 ,
32 ,
1  ,
4  ,
42 ,
53 ,
24 ,
26 ,
44 ,
58 ,
24 ,
33 ,
32 ,
22 ,
28 ,
5  ,
21 ,
13 ,
53 ,
83 ,
43 ,
14 ,
4  ,
26 ,
36 ,
25 ,
61 ,
34 ,
12 ,
61 ,
34 ,
23 ,
14 ,
25 ,
31 ,
26 ,
22 ,
42 ,
41 ,
27 ,
35 ,
56 ,
75 ,
15 ,
87 ,
33 ,
12 ,
4  ,
7  ,
15 ,
35 ,
53 ,
14 ,
45 ,
22 ,
16 ,
4  ,
36 ,
34 ,
5  ,
27 ,
24 ,
26 ,
46 ,
38 ,
43 ,
12 ,
23 ,
55 ,
24 ,
25 ,
36 ,
47 ,
17 ,
46 ,
16 ,
28 ,
34 ,
27 ,
37 ,
15 ,
35 ,
5  ,
18 ,
43 ,
76 ,
45 ,
32 ,
48 ,
26 ,
47 ,
57 ,
37 ,
58 ,
25 ,
28 ,
36 ,
16 ,
17 ,
18 ,
29 ,
5  ,
45 ,
35 ,
6  ,
46 ,
38 ,
40 ,
19 ,
27 ,
18 ,
38 ,
8  ,
48 ,
29 ,
26 ,
19 ,
39 ,
9  ,
30 ,
6  ,
14 ,
49 ,
45 ,
68 ,
70 ,
58 ,
40 ,
17 ,
39 ,
24 ,
19 ,
30 ,
20 ,
10 ,
28 ,
68 ,
26 ,
58 ,
27 ,
38 ,
50 ,
49 ,
37 ,
60 ,
35 ,
59 ,
40 ,
9  ,
29 ,
40 ,
20 ,
28 ,
50 ,
60 ,
59 ,
38 ,
39 ,
10 ,
18 ,
27 ,
9  ,
68 ,
80 ,
19 ,
26 ,
17 ,
47 ,
48 ,
22 ,
51 ,
42 ,
11 ,
21 ,
41 ,
61 ,
33 ,
53 ,
32 ,
23 ,
34 ,
83 ,
2  ,
1  ,
12 ,
43 ,
62 ,
63 ,
35 ,
34 ,
31 ,
42 ,
22 ,
43 ,
5  ,
41 ,
21 ,
64 ,
44 ,
52 ,
33 ,
63 ,
14 ,
51 ,
12 ,
13 ,
23 ,
36 ,
15 ,
43 ,
32 ,
13 ,
34 ,
52 ,
23 ,
22 ,
31 ,
53 ,
35 ,
71 ,
24 ,
46 ,
20 ,
44 ,
42 ,
25 ,
45 ,
64 ,
21 ,
35 ,
33 ,
38 ,
54 ,
24 ,
53 ,
44 ,
31 ,
14 ,
74 ,
56 ,
23 ,
37 ,
27 ,
45 ,
25 ,
62 ,
43 ,
42 ,
65 ,
25 ,
45 ,
57 ,
36 ,
24 ,
38 ,
56 ,
34 ,
22 ,
28 ,
47 ,
37 ,
55 ,
31 ,
21 ,
33 ,
41 ,
14 ,
76 ,
48 ,
26 ,
46 ,
37 ,
38 ,
35 ,
15 ,
16 ,
27 ,
56 ,
34 ,
25 ,
47 ,
39 ,
24 ,
32 ,
33 ,
7  ,
43 ,
23 ,
6  ,
36 ,
27 ,
47 ,
56 ,
26 ,
38 ,
46 ,
15 ,
39 ,
17 ,
77 ,
35 ,
58 ,
48 ,
28 ,
57 ,
18 ,
34 ,
23 ,
45 ,
68 ,
59 ,
49 ,
8  ,
37 ,
40 ,
28 ,
29 ,
27 ,
18 ,
48 ,
36 ,
39 ,
70 ,
17 ,
7  ,
6  ,
47 ,
25 ,
78 ,
48 ,
29 ,
49 ,
50 ,
40 ,
38 ,
28 ,
57 ,
16 ,
9  ,
58 ,
59 ,
27 ,
37 ,
19 ,
26 ,
80 ,
30 ,
60 ,
20 ,
50 ,
20 ,
39 ,
30 ,
38 ,
19 ,
29 ,
90 ,
26 ,
49 ,
60 ,
76 ,
70 ,
48 ,
10 ,
28 ,
57 ,
47 ,
59 ,
89 ,
42 ,
43 ,
31 ,
33 ,
62 ,
51 ,
22 ,
32 ,
61 ,
52 ,
21 ,
71 ,
53 ,
11 ,
63 ,
73 ,
2  ,
44 ,
16 ,
45 ,
52 ,
41 ,
53 ,
63 ,
43 ,
62 ,
32 ,
44 ,
21 ,
31 ,
51 ,
61 ,
22 ,
33 ,
81 ,
71 ,
72 ,
55 ,
12 ,
83 ,
33 ,
53 ,
42 ,
3  ,
34 ,
13 ,
14 ,
32 ,
64 ,
41 ,
62 ,
44 ,
31 ,
85 ,
73 ,
12 ,
22 ,
24 ,
63 ,
54 ,
34 ,
83 ,
24 ,
42 ,
54 ,
66 ,
41 ,
43 ,
56 ,
55 ,
68 ,
84 ,
64 ,
45 ,
46 ,
33 ,
53 ,
12 ,
74 ,
63 ,
55 ,
95 ,
23 ,
78 ,
35 ,
44 ,
65 ,
43 ,
42 ,
46 ,
63 ,
25 ,
56 ,
48 ,
36 ,
47 ,
85 ,
33 ,
57 ,
54 ,
37 ,
89 ,
45 ,
56 ,
38 ,
47 ,
66 ,
36 ,
26 ,
35 ,
69 ,
24 ,
48 ,
67 ,
44 ,
55 ,
43 ,
17 ,
77 ,
49 ,
77 ,
27 ,
56 ,
49 ,
68 ,
39 ,
55 ,
57 ,
16 ,
44 ,
17 ,
37 ,
48 ,
65 ,
59 ,
36 ,
46 ,
45 ,
7  ,
67 ,
39 ,
49 ,
58 ,
47 ,
60 ,
28 ,
68 ,
38 ,
27 ,
59 ,
50 ,
37 ,
78 ,
26 ,
40 ,
55 ,
66 ,
69 ,
57 ,
67 ,
50 ,
70 ,
39 ,
38 ,
58 ,
59 ,
36 ,
48 ,
57 ,
69 ,
30 ,
78 ,
29 ,
99 ,
47 ,
18 ,
46 ,
19 ,
67 ,
68 ,
49 ,
30 ,
40 ,
87 ,
65 ,
60 ,
48 ,
59 ,
78 ,
70 ,
39 ,
47 ,
57 ,
46 ,
36 ,
19 ,
8  ,
25 ,
69 ,
80 ,
52 ,
61 ,
41 ,
71 ,
81 ,
21 ,
62 ,
42 ,
31 ,
12 ,
63 ,
57 ,
82 ,
83 ,
35 ,
72 ,
43 ,
46 ,
53 ,
54 ,
53 ,
42 ,
62 ,
32 ,
54 ,
61 ,
72 ,
51 ,
41 ,
71 ,
63 ,
64 ,
66 ,
55 ,
34 ,
31 ,
73 ,
46 ,
65 ,
81 ,
52 ,
55 ,
45 ,
64 ,
73 ,
41 ,
54 ,
63 ,
43 ,
97 ,
72 ,
62 ,
51 ,
81 ,
33 ,
22 ,
23 ,
3  ,
67 ,
12 ,
44 ,
45 ,
64 ,
62 ,
55 ,
67 ,
53 ,
51 ,
52 ,
42 ,
43 ,
12 ,
58 ,
74 ,
76 ,
56 ,
63 ,
68 ,
72 ,
24 ,
57 ,
67 ,
37 ,
53 ,
65 ,
35 ,
22 ,
45 ,
54 ,
56 ,
24 ,
74 ,
75 ,
40 ,
52 ,
47 ,
25 ,
73 ,
43 ,
34 ,
57 ,
27 ,
55 ,
66 ,
65 ,
46 ,
54 ,
58 ,
43 ,
77 ,
16 ,
26 ,
68 ,
87 ,
44 ,
36 ,
47 ,
76 ,
53 ,
86 ,
46 ,
47 ,
56 ,
67 ,
87 ,
66 ,
37 ,
79 ,
58 ,
59 ,
55 ,
86 ,
35 ,
68 ,
65 ,
48 ,
27 ,
26 ,
54 ,
45 ,
57 ,
38 ,
47 ,
60 ,
30 ,
46 ,
59 ,
40 ,
78 ,
56 ,
68 ,
20 ,
85 ,
49 ,
69 ,
28 ,
48 ,
87 ,
17 ,
77 ,
69 ,
57 ,
60 ,
39 ,
49 ,
99 ,
58 ,
80 ,
56 ,
70 ,
98 ,
29 ,
40 ,
68 ,
48 ,
88 ,
55 ,
50 ,
90 ,
28 ,
49 ,
70 ,
79 ,
59 ,
47 ,
68 ,
39 ,
58 ,
50 ,
48 ,
69 ,
56 ,
28 ,
30 ,
80 ,
67 ,
40 ,
66 ,
78 ,
88 ,
51 ,
73 ,
62 ,
71 ,
81 ,
53 ,
52 ,
92 ,
31 ,
41 ,
82 ,
72 ,
63 ,
74 ,
42 ,
91 ,
85 ,
83 ,
23 ,
64 ,
61 ,
72 ,
63 ,
82 ,
64 ,
91 ,
73 ,
52 ,
74 ,
45 ,
25 ,
42 ,
53 ,
32 ,
51 ,
92 ,
71 ,
55 ,
75 ,
43 ,
65 ,
62 ,
72 ,
44 ,
43 ,
74 ,
61 ,
64 ,
83 ,
73 ,
71 ,
53 ,
67 ,
93 ,
57 ,
82 ,
84 ,
95 ,
55 ,
81 ,
63 ,
84 ,
65 ,
53 ,
92 ,
93 ,
74 ,
34 ,
66 ,
54 ,
94 ,
73 ,
43 ,
78 ,
55 ,
67 ,
77 ,
68 ,
51 ,
45 ,
73 ,
64 ,
66 ,
85 ,
55 ,
75 ,
33 ,
67 ,
83 ,
44 ,
86 ,
46 ,
76 ,
45 ,
87 ,
63 ,
57 ,
54 ,
47 ,
53 ,
76 ,
34 ,
67 ,
65 ,
15 ,
77 ,
46 ,
56 ,
59 ,
75 ,
86 ,
55 ,
85 ,
74 ,
64 ,
89 ,
21 ,
72 ,
57 ,
63 ,
77 ,
53 ,
76 ,
97 ,
66 ,
47 ,
46 ,
55 ,
57 ,
69 ,
68 ,
64 ,
27 ,
58 ,
49 ,
65 ,
87 ,
59 ,
78 ,
89 ,
77 ,
67 ,
58 ,
76 ,
60 ,
59 ,
78 ,
57 ,
69 ,
47 ,
88 ,
79 ,
70 ,
97 ,
99 ,
65 ,
74 ,
98 ,
48 ,
66 ,
68 ,
80 ,
70 ,
59 ,
79 ,
89 ,
50 ,
60 ,
67 ,
48 ,
78 ,
49 ,
65 ,
37 ,
57 ,
38 ,
58 ,
56 ,
98 ,
20 ,
49 ,
66 ,
60 ,
100,
69 ,
59 ,
85 ,
80 ,
77 ,
50 ,
20 ,
78 ,
79 ,
90 ,
67 ,
30 ,
68 ,
88 ,
99 ,
58 ,
72 ,
81 ,
85 ,
74 ,
82 ,
73 ,
91 ,
62 ,
42 ,
63 ,
61 ,
67 ,
51 ,
43 ,
92 ,
83 ,
41 ,
52 ,
93 ,
31 ,
62 ,
71 ,
52 ,
24 ,
73 ,
81 ,
82 ,
61 ,
47 ,
63 ,
51 ,
42 ,
83 ,
75 ,
45 ,
53 ,
91 ,
33 ,
46 ,
74 ,
72 ,
63 ,
74 ,
54 ,
52 ,
93 ,
83 ,
75 ,
62 ,
85 ,
82 ,
64 ,
71 ,
44 ,
56 ,
84 ,
43 ,
81 ,
53 ,
94 ,
84 ,
65 ,
54 ,
73 ,
76 ,
75 ,
94 ,
85 ,
72 ,
48 ,
83 ,
62 ,
64 ,
63 ,
77 ,
98 ,
34 ,
71 ,
82 ,
44 ,
65 ,
55 ,
85 ,
86 ,
74 ,
44 ,
96 ,
73 ,
84 ,
95 ,
77 ,
76 ,
94 ,
62 ,
97 ,
66 ,
99 ,
54 ,
57 ,
56 ,
66 ,
78 ,
75 ,
87 ,
99 ,
86 ,
77 ,
39 ,
74 ,
54 ,
95 ,
85 ,
47 ,
35 ,
23 ,
64 ,
55 ,
82 ,
56 ,
80 ,
76 ,
78 ,
69 ,
67 ,
66 ,
59 ,
95 ,
68 ,
35 ,
74 ,
88 ,
97 ,
58 ,
57 ,
27 ,
98 ,
79 ,
87 ,
96 ,
80 ,
58 ,
79 ,
77 ,
88 ,
74 ,
76 ,
48 ,
90 ,
80 ,
14 ,
98 ,
68 ,
69 ,
67 ,
87 ,
97 ,
35 ,
70 ,
89 ,
66 ,
97 ,
68 ,
78 ,
99 ,
80 ,
100,
98 ,
60 ,
67 ,
76 ,
89 ,
69 ,
59 ,
70 ,
30 ,
77 ,
88 ,
75 ,
49 ,
58 ,
60 ,
100,
79 ,
70 ,
68 ,
89 ,
88 ,
48 ,
90 ,
77 ,
69 ,
78 ,
76 ,
75 ,
86 ,
59 ,
27 ,
98 ,
12 ,
20 ,
71 ,
91 ,
92 ,
82 ,
93 ,
61 ,
63 ,
51 ,
53 ,
42 ,
73 ,
52 ,
83 ,
43 ,
72 ,
84 ,
74 ,
96 ,
44 ,
54 ,
92 ,
85 ,
72 ,
83 ,
62 ,
52 ,
81 ,
34 ,
94 ,
84 ,
93 ,
73 ,
91 ,
74 ,
63 ,
71 ,
61 ,
86 ,
53 ,
42 ,
84 ,
53 ,
74 ,
94 ,
82 ,
93 ,
72 ,
92 ,
63 ,
52 ,
85 ,
73 ,
87 ,
65 ,
81 ,
61 ,
43 ,
62 ,
95 ,
98 ,
82 ,
83 ,
64 ,
93 ,
75 ,
74 ,
94 ,
85 ,
96 ,
95 ,
86 ,
54 ,
65 ,
73 ,
76 ,
62 ,
55 ,
72 ,
67 ,
63 ,
96 ,
84 ,
92 ,
63 ,
56 ,
95 ,
86 ,
55 ,
76 ,
74 ,
88 ,
83 ,
75 ,
94 ,
77 ,
67 ,
62 ,
65 ,
64 ,
97 ,
96 ,
76 ,
87 ,
66 ,
88 ,
95 ,
85 ,
97 ,
77 ,
68 ,
90 ,
57 ,
75 ,
28 ,
74 ,
84 ,
98 ,
45 ,
93 ,
56 ,
88 ,
91 ,
77 ,
96 ,
76 ,
86 ,
68 ,
89 ,
85 ,
97 ,
98 ,
99 ,
79 ,
67 ,
69 ,
90 ,
75 ,
47 ,
78 ,
84 ,
90 ,
98 ,
78 ,
87 ,
68 ,
99 ,
86 ,
94 ,
66 ,
59 ,
89 ,
69 ,
100,
85 ,
97 ,
67 ,
70 ,
84 ,
65 ,
80 ,
79 ,
90 ,
87 ,
88 ,
99 ,
97 ,
100,
78 ,
69 ,
59 ,
76 ,
68 ,
80 ,
77 ,
58 ,
66 ,
98 ,
67 ,
96 ,
86 ,
79 ,
100,
89 ,
80 ,
88 ,
76 ,
87 ,
99 ,
66 ,
68 ,
58 ,
70 ,
69 ,
78 ,
86 ,
60 ,
59 ,
98 ,
77 ,
97 ,
82 ,
71 ,
92 ,
81 ,
64 ,
93 ,
84 ,
72 ,
94 ,
83 ,
63 ,
73 ,
62 ,
96 ,
61 ,
95 ,
52 ,
74 ,
51 ,
53 ,
93 ,
91 ,
82 ,
83 ,
84 ,
55 ,
94 ,
71 ,
95 ,
86 ,
52 ,
44 ,
73 ,
64 ,
72 ,
81 ,
63 ,
61 ,
62 ,
85 ,
81 ,
82 ,
92 ,
83 ,
97 ,
94 ,
73 ,
65 ,
91 ,
72 ,
84 ,
85 ,
95 ,
75 ,
98 ,
53 ,
88 ,
74 ,
96 ,
63 ,
73 ,
84 ,
74 ,
93 ,
95 ,
96 ,
75 ,
85 ,
62 ,
97 ,
92 ,
72 ,
81 ,
83 ,
64 ,
99 ,
82 ,
54 ,
91 ,
87 ,
85 ,
96 ,
84 ,
92 ,
88 ,
94 ,
86 ,
97 ,
75 ,
77 ,
81 ,
93 ,
99 ,
74 ,
65 ,
83 ,
71 ,
87 ,
56 ,
55 ,
97 ,
86 ,
94 ,
54 ,
75 ,
95 ,
76 ,
74 ,
98 ,
85 ,
87 ,
65 ,
56 ,
66 ,
78 ,
57 ,
88 ,
37 ,
83 ,
99 ,
88 ,
85 ,
96 ,
98 ,
78 ,
77 ,
95 ,
58 ,
99 ,
87 ,
86 ,
90 ,
92 ,
89 ,
67 ,
94 ,
68 ,
60 ,
76 ,
75 ,
99 ,
87 ,
78 ,
89 ,
100,
96 ,
97 ,
95 ,
86 ,
68 ,
88 ,
80 ,
70 ,
77 ,
79 ,
74 ,
57 ,
90 ,
66 ,
69 ,
89 ,
100,
98 ,
88 ,
68 ,
79 ,
97 ,
87 ,
67 ,
90 ,
69 ,
80 ,
95 ,
78 ,
59 ,
77 ,
96 ,
50 ,
76 ,
85 ,
99 ,
98 ,
90 ,
80 ,
79 ,
89 ,
70 ,
69 ,
76 ,
78 ,
88 ,
59 ,
84 ,
87 ,
97 ,
95 ,
94 ,
77 ,
60 ,
39 );

end package wm_package; 
package body wm_package is
 
  
end package body wm_package;
